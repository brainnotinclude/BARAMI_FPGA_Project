`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/12 18:29:06
// Design Name: 
// Module Name: gfx
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module gfx(
    input wire [11:0] i_x,
    input wire [11:0] i_y,
    input wire pix_clk,
    input wire [6:0] character,
    
    output wire [7:0] o_red,
    output wire [7:0] o_blue,
    output wire [7:0] o_green
    );
    
    reg pixval;
    wire [3:0] res_x;
    wire [3:0] res_y;
    
    localparam [0:15][0:15] zero = {
   //0 => you can draw 1, ...,9, +, -, *, /, % like this
       4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,
       4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
   };
   
    localparam [0:15][0:15] one = {

4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0

        
   };

    localparam [0:15][0:15] two = {
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd1,	4'd0,	4'd0,
4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0,	4'd0
   };
    localparam [0:15][0:15] three = {
       
   };
    localparam [0:15][0:15] four = {
       
   };
    localparam [0:15][0:15] five = {
       
   };
    localparam [0:15][0:15] six = {
       
   };
    localparam [0:15][0:15] seven = {
       
   };
    localparam [0:15][0:15] eight = {
       
   };
    localparam [0:15][0:15] nine = {
       
   };
    localparam [0:15][0:15] plus = {
       
   };
    localparam [0:15][0:15] minus = {
       
   };
    localparam [0:15][0:15] product = {
       
   };
    localparam [0:15][0:15] divide = {
       
   };
    localparam [0:15][0:15] modular = {
       
   };
    localparam [0:15][0:15] equalSign = {
       
   };
   
   assign res_x = i_x%16;
   assign res_y = i_y%16;
   
   always@(*) begin
       case(character)
           7'h30: pixval = zero[res_x][res_y];
           7'h31: pixval = one[res_x][res_y];
           7'h32: pixval = two[res_x][res_y];
           7'h33: pixval = three[res_x][res_y];
           7'h34: pixval = four[res_x][res_y];
           7'h35: pixval = five[res_x][res_y];
           7'h36: pixval = six[res_x][res_y];
           7'h37: pixval = seven[res_x][res_y];
           7'h38: pixval = eight[res_x][res_y];
           7'h39: pixval = nine[res_x][res_y];
           7'h2B: pixval = plus[res_x][res_y];
           7'h2D: pixval = minus[res_x][res_y];
           7'h2A: pixval = product[res_x][res_y];
           7'h2F: pixval = divide[res_x][res_y];
           7'h25: pixval = modular[res_x][res_y];
           default: pixval = 1'b0;                      //Black
       endcase
   end
   
   //white if 1, black if 0
   assign o_red = pixval ? 8'hFF: 8'h00;
   assign o_green = pixval ? 8'hFF: 8'h00;
   assign o_blue = pixval ? 8'hFF: 8'h00;
    
endmodule
